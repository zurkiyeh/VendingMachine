library verilog;
use verilog.vl_types.all;
entity Vending_Machine_vlg_vec_tst is
end Vending_Machine_vlg_vec_tst;
